module types

pub struct ErrorMsg {
	msg  string
	code int
}
