module main

pub fn on_panic() {
	print_backtrace()
}
