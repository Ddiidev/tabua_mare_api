module web_ctx

import veb

pub struct WebCtx {
	veb.Context
}
