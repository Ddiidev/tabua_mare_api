module web_ctx

import veb

pub struct WsCtx {
	veb.Context
}
