module dto

pub struct DTOHaborMareListHaborNameByState {
pub:
	id                          int    @[omitempty]
	year                        int    @[omitempty]
	harbor_name                 string @[omitempty]
	data_collection_institution string @[omitempty]
}
