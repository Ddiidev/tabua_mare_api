module constants

import time

pub const year = time.now().year
