module types

pub type UUID = string
