module auth_user

// UserData representa os dados do usuário para o JWT
pub struct UserData {
pub:
	email string
	name  string
}
