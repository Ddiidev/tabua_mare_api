module components_view

pub struct ComponentsView {}
